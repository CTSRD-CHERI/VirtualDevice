/*-
 * Copyright (c) 2022 Jonathan Woodruff
 * All rights reserved.
 *
 * @BERiLICENSE_HEADER_START@
 *
 * Licensed to BERI Open Systems C.I.C. (BERI) under one or more contributor
 * license agreements.  See the NOTICE file distributed with this work for
 * additional information regarding copyright ownership.  BERI licenses this
 * file to you under the BERI Hardware-Software License, Version 1.0 (the
 * "License"); you may not use this file except in compliance with the
 * License.  You may obtain a copy of the License at:
 *
 *   http://www.beri-open-systems.org/legal/license-1-0.txt
 *
 * Unless required by applicable law or agreed to in writing, Work distributed
 * under the License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied.  See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * @BERiLICENSE_HEADER_END@
 */
 
import VirtualDevice::*;
import AXI4::*;
import SourceSink::*;
 
(*synthesize*)
module mkTestVirtualDevice();
  VirtualDeviceIfc#(2,32,64) vd <- mkVirtualDevice;
  
  rule virtualRequest;
    AXI4_ARFlit#(2,32,0) readFlit = defaultValue;
    readFlit.araddr = 0;
    vd.virt.ar.put(readFlit);
    $display("Put one in virt: ", fshow(readFlit));
  endrule
  
  rule virtualResponse(vd.virt.r.canPeek);
    $display("Look at me! ", fshow(vd.virt.r.peek));
    vd.virt.r.drop;
  endrule
  
  rule managementRequest;
  endrule
  
  rule managementResponse;
  endrule
endmodule
